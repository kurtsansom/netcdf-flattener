netcdf input4 {

// global attributes:
		:Conventions = "CF-1.8" ;

group: group1 {
  dimensions:
  	lat = 5 ;
  	bounds2 = 2 ;
  	lon = 8 ;
  variables:
  	double lat_bnds(lat, bounds2) ;
  	double lat(lat) ;
  		lat:units = "degrees_north" ;
  		lat:standard_name = "latitude" ;
  		lat:bounds = "lat_bnds" ;
  	double lon_bnds(lon, bounds2) ;
  	double lon(lon) ;
  		lon:units = "degrees_east" ;
  		lon:standard_name = "longitude" ;
  		lon:bounds = "lon_bnds" ;
  	double time ;
  		time:units = "days since 2018-12-01" ;
  		time:standard_name = "time" ;
  	double q(lat, lon) ;
  		q:project = "research" ;
  		q:standard_name = "specific_humidity" ;
  		q:units = "1" ;
  		q:coordinates = "time" ;
  		q:cell_methods = "area: mean any_valid_name: mean time: mean bounds2: mean" ;
  data:

   lat_bnds =
  -90, -60,
  -60, -30,
  -30, 30,
  30, 60,
  60, 90 ;

   lat = -75, -45, 0, 45, 75 ;

   lon_bnds =
  0, 45,
  45, 90,
  90, 135,
  135, 180,
  180, 225,
  225, 270,
  270, 315,
  315, 360 ;

   lon = 22.5, 67.5, 112.5, 157.5, 202.5, 247.5, 292.5, 337.5 ;

   time = 31 ;

   q =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013 ;
  } // group group1
}
