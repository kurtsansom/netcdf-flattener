// -*-C++-*-
// Generate netCDF file with:
// ncgen -k netCDF-4 -b -o ~/nco/data/cf_grp.nc ~/nco/data/cf

netcdf input1 {
dimensions:
	lat = 180 ;
	lon = 360 ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:title = "A template/test dataset for Groups in CF" ;
		:history = "Global history attribute" ;

group: e3sm {
  dimensions:
  	lat = 2 ;
  	lon = 3 ;
  	time = UNLIMITED ; // (4 currently)
  variables:
  	double lat(lat) ;
  		lat:long_name = "latitude" ;
  		lat:standard_name = "latitude" ;
  		lat:units = "degrees_north" ;
  		lat:axis = "Y" ;
  	double lon(lon) ;
  		lon:long_name = "longitude" ;
  		lon:standard_name = "longitude" ;
  		lon:units = "degrees_east" ;
  		lon:axis = "X" ;
  	double time(time) ;
  		time:long_name = "time of measurement" ;
  		time:standard_name = "time" ;
  		time:units = "days since 1964-03-12 12:09:00 -9:00" ;
  		time:calendar = "leap" ;

  // group attributes:
  		:title = "group-level title attribute is allowed" ;
  data:

   lat = -90, 90 ;

   lon = 0, 120, 240 ;

   time = 1, 2, 3, 4 ;

  group: e3sm_01 {
    variables:
    	float tas(time, lat, lon) ;
    		tas:long_name = "surface air temperature" ;
    		tas:standard_name = "air_temperature" ;
    		tas:units = "kelvin" ;
    		tas:coordinates = "time lat lon" ;

    // group attributes:
    		:Realization = "1" ;
    		:history = "Group-level history attributes are OK too" ;
    data:

     tas =
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15 ;
    } // group e3sm_01

  group: e3sm_02 {
    variables:
    	float tas(time, lat, lon) ;
    		tas:long_name = "surface air temperature" ;
    		tas:standard_name = "air_temperature" ;
    		tas:coordinates = "/e3sm/time /e3sm/lat /e3sm/lon" ;

    // group attributes:
    		:Realization = "2" ;
    data:

     tas =
  272.15, 272.15, 272.15,
  272.15, 272.15, 272.15,
  272.15, 272.15, 272.15,
  272.15, 272.15, 272.15,
  272.15, 272.15, 272.15,
  272.15, 272.15, 272.15,
  272.15, 272.15, 272.15,
  272.15, 272.15, 272.15 ;
    } // group e3sm_02

  group: e3sm_03 {
    variables:
    	float tas(time, lat, lon) ;
    		tas:long_name = "surface air temperature" ;
    		tas:standard_name = "air_temperature" ;
    		tas:coordinates = "../time ../lat ../lon" ;

    // group attributes:
    		:Realization = "3" ;
    data:

     tas =
  273.15, 273.15, 273.15,
  273.15, 273.15, 273.15,
  273.15, 273.15, 273.15,
  273.15, 273.15, 273.15,
  273.15, 273.15, 273.15,
  273.15, 273.15, 273.15,
  273.15, 273.15, 273.15,
  273.15, 273.15, 273.15 ;
    } // group e3sm_03
  } // group e3sm

group: nasa {
  dimensions:
  	lat = 2 ;
  	lon = 3 ;
  	time = UNLIMITED ; // (4 currently)

  group: nasa_data {
    variables:
    	float tas(time, lat, lon) ;
    		tas:long_name = "surface air temperature" ;
    		tas:standard_name = "air_temperature" ;
    		tas:units = "kelvin" ;
    		tas:coordinates = "time lat lon" ;
    	float sic(time, lat, lon) ;
    		sic:long_name = "sea-ice concentration" ;
    		sic:standard_name = "sea_ice_area_fraction" ;
    		sic:units = "1" ;
    		sic:coordinates = "/nasa/nasa_geo/time /nasa/nasa_geo/lat /nasa/nasa_geo/lon" ;
    	float sit(time, lat, lon) ;
    		sit:long_name = "sea-ice thickness" ;
    		sit:standard_name = "sea_ice_thickness" ;
    		sit:units = "meter" ;
    		sit:coordinates = "../nasa_geo/time ../nasa_geo/lat ../nasa_geo/lon" ;

    // group attributes:
    		:history = "Group-level history attributes are OK too" ;
    data:

     tas =
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15 ;

     sic =
  0.73, 0.73, 0.73,
  0.73, 0.73, 0.73,
  0.73, 0.73, 0.73,
  0.73, 0.73, 0.73,
  0.73, 0.73, 0.73,
  0.73, 0.73, 0.73,
  0.73, 0.73, 0.73,
  0.73, 0.73, 0.73 ;

     sit =
  3.7, 3.7, 3.7,
  3.7, 3.7, 3.7,
  3.7, 3.7, 3.7,
  3.7, 3.7, 3.7,
  3.7, 3.7, 3.7,
  3.7, 3.7, 3.7,
  3.7, 3.7, 3.7,
  3.7, 3.7, 3.7 ;
    } // group nasa_data

  group: nasa_geo {
    variables:
    	double lat(lat) ;
    		lat:long_name = "latitude" ;
    		lat:standard_name = "latitude" ;
    		lat:units = "degrees_north" ;
    		lat:axis = "Y" ;
    	double lon(lon) ;
    		lon:long_name = "longitude" ;
    		lon:standard_name = "longitude" ;
    		lon:units = "degrees_east" ;
    		lon:axis = "X" ;
    	double time(time) ;
    		time:long_name = "time of measurement" ;
    		time:standard_name = "time" ;
    		time:units = "days since 1964-03-12 12:09:00 -9:00" ;
    		time:calendar = "leap" ;
    data:

     lat = -90, 90 ;

     lon = 0, 120, 240 ;

     time = 1, 2, 3, 4 ;
    } // group nasa_geo
  } // group nasa

group: nsidc {
  dimensions:
  	time = UNLIMITED ; // (5 currently)

  group: nsidc {
    variables:
    	float tas(time) ;
    		tas:long_name = "surface air temperature" ;
    		tas:standard_name = "air_temperature" ;
    		tas:units = "kelvin" ;
    	double time(time) ;
    		time:long_name = "time of measurement" ;
    		time:standard_name = "time" ;
    		time:units = "days since 1964-03-12 12:09:00 -9:00" ;
    		time:calendar = "leap" ;
    data:

     tas = 274.15, 274.15, 274.15, 274.15, 274.15 ;

     time = 1, 2, 3, 4, 5 ;
    } // group nsidc
  } // group nsidc
}
