netcdf output2 {

// global attributes:
                :group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890\#group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890\#attr_short_234567890123456789012345678901234567890123 = "This attribute name would be flattened as 255 character long." ;
                :\6976e5b3f72cd92fa88d106c519b9739c399ef89\#attr_exact_2345678901234567890123456789012345678901234 = "This attribute name would be flattened as 256 character long." ;
                :\6976e5b3f72cd92fa88d106c519b9739c399ef89\#attr_long1_23456789012345678901234567890123456789012345 = "This attribute name would be flattened as 257 character long." ;
                :\6976e5b3f72cd92fa88d106c519b9739c399ef89\#attr_long2_23456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234 = "This attribute name would be flattened as 416 character long, and with hashing the path would be 255 characters long." ;
                :ebeb0ce7276e1c4a5d72e6f4ba20b0e96f992b3b = "This attribute name would be flattened as 417 characters long, and with hashing the path would be 256 characters long." ;
                string :flattener_name_mapping_attributes = "group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890#group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890#attr_short_234567890123456789012345678901234567890123: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_short_234567890123456789012345678901234567890123", "6976e5b3f72cd92fa88d106c519b9739c399ef89#attr_exact_2345678901234567890123456789012345678901234: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_exact_2345678901234567890123456789012345678901234", "6976e5b3f72cd92fa88d106c519b9739c399ef89#attr_long1_23456789012345678901234567890123456789012345: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_long1_23456789012345678901234567890123456789012345", "6976e5b3f72cd92fa88d106c519b9739c399ef89#attr_long2_23456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_long2_23456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234", "ebeb0ce7276e1c4a5d72e6f4ba20b0e96f992b3b: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_long3_234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345" ;
                :flattener_name_mapping_dimensions = "" ;
                :flattener_name_mapping_variables = "" ;
                :_NCProperties = "version=2,netcdf=4.6.3,hdf5=1.10.4" ;
}
