netcdf output4 {
dimensions:
	group1\#lat = 5 ;
	group1\#bounds2 = 2 ;
	group1\#lon = 8 ;
variables:
	double group1\#lat_bnds(group1\#lat, group1\#bounds2) ;
	double group1\#lat(group1\#lat) ;
		group1\#lat:units = "degrees_north" ;
		group1\#lat:standard_name = "latitude" ;
		group1\#lat:bounds = "group1#lat_bnds" ;
	double group1\#lon_bnds(group1\#lon, group1\#bounds2) ;
	double group1\#lon(group1\#lon) ;
		group1\#lon:units = "degrees_east" ;
		group1\#lon:standard_name = "longitude" ;
		group1\#lon:bounds = "group1#lon_bnds" ;
	double group1\#time ;
		group1\#time:units = "days since 2018-12-01" ;
		group1\#time:standard_name = "time" ;
	double group1\#q(group1\#lat, group1\#lon) ;
		group1\#q:project = "research" ;
		group1\#q:standard_name = "specific_humidity" ;
		group1\#q:units = "1" ;
		group1\#q:coordinates = "group1#time" ;
		group1\#q:cell_methods = "area: mean any_valid_name: mean group1#time: mean group1#bounds2: mean" ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:flattener_name_mapping_attributes = "Conventions: /Conventions" ;
		string :flattener_name_mapping_dimensions = "group1#lat: /group1/lat", "group1#bounds2: /group1/bounds2", "group1#lon: /group1/lon" ;
		string :flattener_name_mapping_variables = "group1#lat_bnds: /group1/lat_bnds", "group1#lat: /group1/lat", "group1#lon_bnds: /group1/lon_bnds", "group1#lon: /group1/lon", "group1#time: /group1/time", "group1#q: /group1/q" ;
data:

 group1\#lat_bnds =
  -90, -60,
  -60, -30,
  -30, 30,
  30, 60,
  60, 90 ;

 group1\#lat = -75, -45, 0, 45, 75 ;

 group1\#lon_bnds =
  0, 45,
  45, 90,
  90, 135,
  135, 180,
  180, 225,
  225, 270,
  270, 315,
  315, 360 ;

 group1\#lon = 22.5, 67.5, 112.5, 157.5, 202.5, 247.5, 292.5, 337.5 ;

 group1\#time = 31 ;

 group1\#q =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013 ;
}
