netcdf output3 {
dimensions:
	lat = 180 ;
	lon = 360 ;
	e3sm\#lat = 2 ;
	e3sm\#lon = 3 ;
	e3sm\#time = UNLIMITED ; // (4 currently)
variables:
	double e3sm\#lat(e3sm\#lat) ;
		e3sm\#lat:long_name = "latitude" ;
		e3sm\#lat:standard_name = "latitude" ;
		e3sm\#lat:units = "degrees_north" ;
		e3sm\#lat:axis = "Y" ;
	double e3sm\#lon(e3sm\#lon) ;
		e3sm\#lon:long_name = "longitude" ;
		e3sm\#lon:standard_name = "longitude" ;
		e3sm\#lon:units = "degrees_east" ;
		e3sm\#lon:axis = "X" ;
	double e3sm\#time(e3sm\#time) ;
		e3sm\#time:long_name = "time of measurement" ;
		e3sm\#time:standard_name = "time" ;
		e3sm\#time:units = "days since 1964-03-12 12:09:00 -9:00" ;
		e3sm\#time:calendar = "leap" ;
	float e3sm\#e3sm_01\#tas(e3sm\#time, e3sm\#lat, e3sm\#lon) ;
		e3sm\#e3sm_01\#tas:long_name = "surface air temperature" ;
		e3sm\#e3sm_01\#tas:standard_name = "air_temperature" ;
		e3sm\#e3sm_01\#tas:units = "kelvin" ;
		e3sm\#e3sm_01\#tas:coordinates = "e3sm#time e3sm#lat e3sm#lon" ;
	float e3sm\#e3sm_01\#sic(e3sm\#time, e3sm\#lat, e3sm\#lon) ;
		e3sm\#e3sm_01\#sic:long_name = "sea-ice concentration" ;
		e3sm\#e3sm_01\#sic:standard_name = "sea_ice_area_fraction" ;
		e3sm\#e3sm_01\#sic:units = "1" ;
		e3sm\#e3sm_01\#sic:coordinates = "e3sm#time REF_NOT_FOUND:_wrong_var e3sm#lon" ;
		e3sm\#e3sm_01\#sic:cell_methods = "REF_NOT_FOUND:_../../../time: mean" ;
		e3sm\#e3sm_01\#sic:cell_measures = "area: REF_NOT_FOUND:_../wrong_group/time" ;
		e3sm\#e3sm_01\#sic:sample_dimension = "REF_NOT_FOUND:_/e3sm/wrong_name" ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:title = "A template/test dataset for Groups in CF" ;
		:history = "Global history attribute" ;
		:e3sm\#title = "group-level title attribute is allowed" ;
		:e3sm\#e3sm_01\#Realization = "1" ;
		:e3sm\#e3sm_01\#history = "Group-level history attributes are OK too" ;
		string :flattener_name_mapping_attributes = "Conventions: /Conventions", "title: /title", "history: /history", "e3sm#title: /e3sm/title", "e3sm#e3sm_01#Realization: /e3sm/e3sm_01/Realization", "e3sm#e3sm_01#history: /e3sm/e3sm_01/history" ;
		string :flattener_name_mapping_dimensions = "lat: /lat", "lon: /lon", "e3sm#lat: /e3sm/lat", "e3sm#lon: /e3sm/lon", "e3sm#time: /e3sm/time" ;
		string :flattener_name_mapping_variables = "e3sm#lat: /e3sm/lat", "e3sm#lon: /e3sm/lon", "e3sm#time: /e3sm/time", "e3sm#e3sm_01#tas: /e3sm/e3sm_01/tas", "e3sm#e3sm_01#sic: /e3sm/e3sm_01/sic" ;
data:

 e3sm\#lat = -90, 90 ;

 e3sm\#lon = 0, 120, 240 ;

 e3sm\#time = 1, 2, 3, 4 ;

 e3sm\#e3sm_01\#tas =
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15 ;

 e3sm\#e3sm_01\#sic =
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15 ;
}
