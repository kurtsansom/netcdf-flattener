netcdf output2 {

// global attributes:
		:group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890__group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890__attr_short_2345678901234567890123456789012345678901 = "This attribute name would be flattened as 255 character long." ;
		:\6976e5b3f72cd92fa88d106c519b9739c399ef89__attr_exact_23456789012345678901234567890123456789012 = "This attribute name would be flattened as 256 character long." ;
		:\6976e5b3f72cd92fa88d106c519b9739c399ef89__attr_long1_234567890123456789012345678901234567890123 = "This attribute name would be flattened as 257 character long." ;
		:\6976e5b3f72cd92fa88d106c519b9739c399ef89__attr_long2_234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012 = "This attribute name would be flattened as 416 character long, and with hashing the path would be 255 characters long." ;
		:aa1dad6fe26a869c57e29e421e6150d7a95235e0 = "This attribute name would be flattened as 417 characters long, and with hashing the path would be 256 characters long." ;
		string :flattener_name_mapping_attributes = "group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890__group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890__attr_short_2345678901234567890123456789012345678901: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_short_2345678901234567890123456789012345678901", "6976e5b3f72cd92fa88d106c519b9739c399ef89__attr_exact_23456789012345678901234567890123456789012: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_exact_23456789012345678901234567890123456789012", "6976e5b3f72cd92fa88d106c519b9739c399ef89__attr_long1_234567890123456789012345678901234567890123: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_long1_234567890123456789012345678901234567890123", "6976e5b3f72cd92fa88d106c519b9739c399ef89__attr_long2_234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_long2_234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012", "aa1dad6fe26a869c57e29e421e6150d7a95235e0: /group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890/attr_long3_23456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234" ;
		:flattener_name_mapping_dimensions = "" ;
		:flattener_name_mapping_variables = "" ;
		:_NCProperties = "version=2,netcdf=4.6.3,hdf5=1.10.4" ;
}
