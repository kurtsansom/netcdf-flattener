netcdf output3 {
dimensions:
	lat = 180 ;
	lon = 360 ;
	e3sm__lat = 2 ;
	e3sm__lon = 3 ;
	e3sm__time = UNLIMITED ; // (4 currently)
variables:
	double e3sm__lat(e3sm__lat) ;
		e3sm__lat:long_name = "latitude" ;
		e3sm__lat:standard_name = "latitude" ;
		e3sm__lat:units = "degrees_north" ;
		e3sm__lat:axis = "Y" ;
	double e3sm__lon(e3sm__lon) ;
		e3sm__lon:long_name = "longitude" ;
		e3sm__lon:standard_name = "longitude" ;
		e3sm__lon:units = "degrees_east" ;
		e3sm__lon:axis = "X" ;
	double e3sm__time(e3sm__time) ;
		e3sm__time:long_name = "time of measurement" ;
		e3sm__time:standard_name = "time" ;
		e3sm__time:units = "days since 1964-03-12 12:09:00 -9:00" ;
		e3sm__time:calendar = "leap" ;
	float e3sm__e3sm_01__tas(e3sm__time, e3sm__lat, e3sm__lon) ;
		e3sm__e3sm_01__tas:long_name = "surface air temperature" ;
		e3sm__e3sm_01__tas:standard_name = "air_temperature" ;
		e3sm__e3sm_01__tas:units = "kelvin" ;
		e3sm__e3sm_01__tas:coordinates = "e3sm__time e3sm__lat e3sm__lon" ;
	float e3sm__e3sm_01__sic(e3sm__time, e3sm__lat, e3sm__lon) ;
		e3sm__e3sm_01__sic:long_name = "sea-ice concentration" ;
		e3sm__e3sm_01__sic:standard_name = "sea_ice_area_fraction" ;
		e3sm__e3sm_01__sic:units = "1" ;
		e3sm__e3sm_01__sic:coordinates = "e3sm__time REF_NOT_FOUND:_wrong_var e3sm__lon" ;
		e3sm__e3sm_01__sic:cell_measures = "area: REF_NOT_FOUND:_../wrong_group/time" ;
		e3sm__e3sm_01__sic:sample_dimension = "REF_NOT_FOUND:_/e3sm/wrong_name" ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:title = "A template/test dataset for Groups in CF" ;
		:history = "Global history attribute" ;
		:e3sm__title = "group-level title attribute is allowed" ;
		:e3sm__e3sm_01__Realization = "1" ;
		:e3sm__e3sm_01__history = "Group-level history attributes are OK too" ;
		string :flattener_name_mapping_attributes = "Conventions: /Conventions", "title: /title", "history: /history", "e3sm__title: /e3sm/title", "e3sm__e3sm_01__Realization: /e3sm/e3sm_01/Realization", "e3sm__e3sm_01__history: /e3sm/e3sm_01/history" ;
		string :flattener_name_mapping_dimensions = "lat: /lat", "lon: /lon", "e3sm__lat: /e3sm/lat", "e3sm__lon: /e3sm/lon", "e3sm__time: /e3sm/time" ;
		string :flattener_name_mapping_variables = "e3sm__lat: /e3sm/lat", "e3sm__lon: /e3sm/lon", "e3sm__time: /e3sm/time", "e3sm__e3sm_01__tas: /e3sm/e3sm_01/tas", "e3sm__e3sm_01__sic: /e3sm/e3sm_01/sic" ;
data:

 e3sm__lat = -90, 90 ;

 e3sm__lon = 0, 120, 240 ;

 e3sm__time = 1, 2, 3, 4 ;

 e3sm__e3sm_01__tas =
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15 ;

 e3sm__e3sm_01__sic =
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15 ;
}
