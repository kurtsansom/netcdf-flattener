// -*-C++-*-
// Generate netCDF file with:
// ncgen -k netCDF-4 -b -o ~/nco/data/cf_grp.nc ~/nco/data/cf

netcdf input3 {
dimensions:
	lat = 180 ;
	lon = 360 ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:title = "A template/test dataset for Groups in CF" ;
		:history = "Global history attribute" ;

group: e3sm {
  dimensions:
  	lat = 2 ;
  	lon = 3 ;
  	time = UNLIMITED ; // (4 currently)
  variables:
  	double lat(lat) ;
  		lat:long_name = "latitude" ;
  		lat:standard_name = "latitude" ;
  		lat:units = "degrees_north" ;
  		lat:axis = "Y" ;
  	double lon(lon) ;
  		lon:long_name = "longitude" ;
  		lon:standard_name = "longitude" ;
  		lon:units = "degrees_east" ;
  		lon:axis = "X" ;
  	double time(time) ;
  		time:long_name = "time of measurement" ;
  		time:standard_name = "time" ;
  		time:units = "days since 1964-03-12 12:09:00 -9:00" ;
  		time:calendar = "leap" ;

  // group attributes:
  		:title = "group-level title attribute is allowed" ;
  data:

   lat = -90, 90 ;

   lon = 0, 120, 240 ;

   time = 1, 2, 3, 4 ;

  group: e3sm_01 {
    variables:
    	float tas(time, lat, lon) ;
    		tas:long_name = "surface air temperature" ;
    		tas:standard_name = "air_temperature" ;
    		tas:units = "kelvin" ;
    		tas:coordinates = "time lat lon" ;
    	float sic(time, lat, lon) ;
    		sic:long_name = "sea-ice concentration" ;
    		sic:standard_name = "sea_ice_area_fraction" ;
    		sic:units = "1" ;
    		sic:coordinates = "time wrong_var lon" ;
    		sic:cell_methods = "../../../time: mean" ;
    		sic:cell_measures = "area: ../wrong_group/time" ;
    		sic:sample_dimension = "/e3sm/wrong_name" ;

    // group attributes:
    		:Realization = "1" ;
    		:history = "Group-level history attributes are OK too" ;
    data:

     tas =
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15 ;
  
     sic =
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15,
  271.15, 271.15, 271.15 ;
    } // group e3sm_01
  } // group e3sm
}
