netcdf output5 {
dimensions:
	group1\#lat = 5 ;
	group1\#lon = 8 ;
	group1\#time = UNLIMITED ; // (6 currently)
variables:
	double group1\#lat(group1\#lat) ;
		group1\#lat:units = "degrees_north" ;
		group1\#lat:standard_name = "latitude" ;
	double group1\#lon(group1\#lon) ;
		group1\#lon:units = "degrees_east" ;
		group1\#lon:standard_name = "longitude" ;
	double group1\#time(group1\#time) ;
		group1\#time:units = "days since 2018-12-01" ;
		group1\#time:standard_name = "time" ;
	double group1\#q1(group1\#time, group1\#lat, group1\#lon) ;
		group1\#q1:standard_name = "specific_humidity" ;
		group1\#q1:units = "1" ;
	double group1\#q2(group1\#time, group1\#lat, group1\#lon) ;
		group1\#q2:standard_name = "specific_humidity" ;
		group1\#q2:units = "1" ;
	double group1\#q3(group1\#time, group1\#lat, group1\#lon) ;
		group1\#q3:standard_name = "specific_humidity" ;
		group1\#q3:units = "1" ;

// global attributes:
		:Conventions = "CF-1.8" ;
		:flattener_name_mapping_attributes = "Conventions: /Conventions" ;
		string :flattener_name_mapping_dimensions = "group1#lat: /group1/lat", "group1#lon: /group1/lon", "group1#time: /group1/time" ;
		string :flattener_name_mapping_variables = "group1#lat: /group1/lat", "group1#lon: /group1/lon", "group1#time: /group1/time", "group1#q1: /group1/q1", "group1#q2: /group1/q2", "group1#q3: /group1/q3" ;
data:

 group1\#lat = -75, -45, 0, 45, 75 ;

 group1\#lon = 22.5, 67.5, 112.5, 157.5, 202.5, 247.5, 292.5, 337.5 ;

 group1\#time = 31, 32, 33, 34, 35, 36 ;

 group1\#q1 =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013,
  1.007, 1.034, 1.003, 1.014, 1.018, 1.037, 1.024, 1.029,
  1.023, 1.036, 1.045, 1.062, 1.046, 1.073, 1.006, 1.066,
  1.11, 1.131, 1.124, 1.146, 1.087, 1.103, 1.057, 1.011,
  1.029, 1.059, 1.039, 1.07, 1.058, 1.072, 1.009, 1.017,
  1.006, 1.036, 1.019, 1.035, 1.018, 1.037, 1.034, 1.013,
  1.007, 1.034, 1.003, 1.014, 1.018, 1.037, 1.024, 1.029,
  1.023, 1.036, 1.045, 1.062, 1.046, 1.073, 1.006, 1.066,
  1.11, 1.131, 1.124, 1.146, 1.087, 1.103, 1.057, 1.011,
  1.029, 1.059, 1.039, 1.07, 1.058, 1.072, 1.009, 1.017,
  1.006, 1.036, 1.019, 1.035, 1.018, 1.037, 1.034, 1.013,
  2.007, 2.034, 2.003, 2.014, 2.018, 2.037, 2.024, 2.029,
  2.023, 2.036, 2.045, 2.062, 2.046, 2.073, 2.006, 2.066,
  2.11, 2.131, 2.124, 2.146, 2.087, 2.103, 2.057, 2.011,
  2.029, 2.059, 2.039, 2.07, 2.058, 2.072, 2.009, 2.017,
  2.006, 2.036, 2.019, 2.035, 2.018, 2.037, 2.034, 2.013,
  3.007, 3.034, 3.003, 3.014, 3.018, 3.037, 3.024, 3.029,
  3.023, 3.036, 3.045, 3.062, 3.046, 3.073, 3.006, 3.066,
  3.11, 3.131, 3.124, 3.146, 3.087, 3.103, 3.057, 3.011,
  3.029, 3.059, 3.039, 3.07, 3.058, 3.072, 3.009, 3.017,
  3.006, 3.036, 3.019, 3.035, 3.018, 3.037, 3.034, 3.013,
  4.007, 4.034, 4.003, 4.014, 4.018, 4.037, 4.024, 4.029,
  4.023, 4.036, 4.045, 4.062, 4.046, 4.073, 4.006, 4.066,
  4.11, 4.131, 4.124, 4.146, 4.087, 4.103, 4.057, 4.011,
  4.029, 4.059, 4.039, 4.07, 4.058, 4.072, 4.009, 4.017,
  4.006, 4.036, 4.019, 4.035, 4.018, 4.037, 4.034, 4.013 ;

 group1\#q2 =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013,
  1.007, 1.034, 1.003, 1.014, 1.018, 1.037, 1.024, 1.029,
  1.023, 1.036, 1.045, 1.062, 1.046, 1.073, 1.006, 1.066,
  1.11, 1.131, 1.124, 1.146, 1.087, 1.103, 1.057, 1.011,
  1.029, 1.059, 1.039, 1.07, 1.058, 1.072, 1.009, 1.017,
  1.006, 1.036, 1.019, 1.035, 1.018, 1.037, 1.034, 1.013,
  1.007, 1.034, 1.003, 1.014, 1.018, 1.037, 1.024, 1.029,
  1.023, 1.036, 1.045, 1.062, 1.046, 1.073, 1.006, 1.066,
  1.11, 1.131, 1.124, 1.146, 1.087, 1.103, 1.057, 1.011,
  1.029, 1.059, 1.039, 1.07, 1.058, 1.072, 1.009, 1.017,
  1.006, 1.036, 1.019, 1.035, 1.018, 1.037, 1.034, 1.013,
  2.007, 2.034, 2.003, 2.014, 2.018, 2.037, 2.024, 2.029,
  2.023, 2.036, 2.045, 2.062, 2.046, 2.073, 2.006, 2.066,
  2.11, 2.131, 2.124, 2.146, 2.087, 2.103, 2.057, 2.011,
  2.029, 2.059, 2.039, 2.07, 2.058, 2.072, 2.009, 2.017,
  2.006, 2.036, 2.019, 2.035, 2.018, 2.037, 2.034, 2.013,
  3.007, 3.034, 3.003, 3.014, 3.018, 3.037, 3.024, 3.029,
  3.023, 3.036, 3.045, 3.062, 3.046, 3.073, 3.006, 3.066,
  3.11, 3.131, 3.124, 3.146, 3.087, 3.103, 3.057, 3.011,
  3.029, 3.059, 3.039, 3.07, 3.058, 3.072, 3.009, 3.017,
  3.006, 3.036, 3.019, 3.035, 3.018, 3.037, 3.034, 3.013,
  4.007, 4.034, 4.003, 4.014, 4.018, 4.037, 4.024, 4.029,
  4.023, 4.036, 4.045, 4.062, 4.046, 4.073, 4.006, 4.066,
  4.11, 4.131, 4.124, 4.146, 4.087, 4.103, 4.057, 4.011,
  4.029, 4.059, 4.039, 4.07, 4.058, 4.072, 4.009, 4.017,
  4.006, 4.036, 4.019, 4.035, 4.018, 4.037, 4.034, 4.013 ;

 group1\#q3 =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013,
  1.007, 1.034, 1.003, 1.014, 1.018, 1.037, 1.024, 1.029,
  1.023, 1.036, 1.045, 1.062, 1.046, 1.073, 1.006, 1.066,
  1.11, 1.131, 1.124, 1.146, 1.087, 1.103, 1.057, 1.011,
  1.029, 1.059, 1.039, 1.07, 1.058, 1.072, 1.009, 1.017,
  1.006, 1.036, 1.019, 1.035, 1.018, 1.037, 1.034, 1.013,
  1.007, 1.034, 1.003, 1.014, 1.018, 1.037, 1.024, 1.029,
  1.023, 1.036, 1.045, 1.062, 1.046, 1.073, 1.006, 1.066,
  1.11, 1.131, 1.124, 1.146, 1.087, 1.103, 1.057, 1.011,
  1.029, 1.059, 1.039, 1.07, 1.058, 1.072, 1.009, 1.017,
  1.006, 1.036, 1.019, 1.035, 1.018, 1.037, 1.034, 1.013,
  2.007, 2.034, 2.003, 2.014, 2.018, 2.037, 2.024, 2.029,
  2.023, 2.036, 2.045, 2.062, 2.046, 2.073, 2.006, 2.066,
  2.11, 2.131, 2.124, 2.146, 2.087, 2.103, 2.057, 2.011,
  2.029, 2.059, 2.039, 2.07, 2.058, 2.072, 2.009, 2.017,
  2.006, 2.036, 2.019, 2.035, 2.018, 2.037, 2.034, 2.013,
  3.007, 3.034, 3.003, 3.014, 3.018, 3.037, 3.024, 3.029,
  3.023, 3.036, 3.045, 3.062, 3.046, 3.073, 3.006, 3.066,
  3.11, 3.131, 3.124, 3.146, 3.087, 3.103, 3.057, 3.011,
  3.029, 3.059, 3.039, 3.07, 3.058, 3.072, 3.009, 3.017,
  3.006, 3.036, 3.019, 3.035, 3.018, 3.037, 3.034, 3.013,
  4.007, 4.034, 4.003, 4.014, 4.018, 4.037, 4.024, 4.029,
  4.023, 4.036, 4.045, 4.062, 4.046, 4.073, 4.006, 4.066,
  4.11, 4.131, 4.124, 4.146, 4.087, 4.103, 4.057, 4.011,
  4.029, 4.059, 4.039, 4.07, 4.058, 4.072, 4.009, 4.017,
  4.006, 4.036, 4.019, 4.035, 4.018, 4.037, 4.034, 4.013 ;
}
